// andEx.v

module andEx( 
		input wire x, y, 
		output wire z
	);

assign z = x & y; // x and y
endmodule