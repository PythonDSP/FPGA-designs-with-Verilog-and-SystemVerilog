// andEx2.v

module andEx2(x, y, z);

input wire x, y;
output wire z;

assign z = x & y;

endmodule 